**********************************************************
* THIS IS nal_nbk_ckt_02_retport.spice for validating the*
* result, which is obtained by the MAPP version.         *   
**********************************************************
r1 1 2 100
r2 1 3 100
r3 2 3 100
r5 3 5 100
r6 4 5 100
r7 4 6 100
r8 5 6 100
*****************
r9 6 7  100k 
r10 6 8 100k
r11 4 7 100k
r12 5 8 100k
r14 7 0 100k
r15 8 0 100k
******************
i13 7 8 dc 0.001
v4 3 4 dc 10
*************************analysis and result**************
.op     
*.tran 0.1m 10m 
*.control
*run 
*plot v(1) 
*.endc 
.end
